`define DW 32	// Data width
`define AW 9	// Address width
`define MD 256	// Memory depth

