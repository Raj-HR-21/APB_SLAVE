
`include "defines.sv"
package apb_slv_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "apb_slv_seq_item.sv"
	`include "apb_slv_sequence.sv"
	`include "apb_slv_sequencer.sv"
	`include "apb_slv_driver.sv"
	`include "apb_slv_monitor.sv"	
	`include "apb_slv_agent.sv"
	`include "apb_slv_scb.sv"
	`include "apb_slv_func_cov.sv"
	`include "apb_slv_environment.sv"
	`include "apb_slv_test.sv"

endpackage
